module AXI2SPI_tb();


endmodule
