module round #(
    parameter DATA_WIDTH = 128;
) (
    input clk;
    input [DATA_WIDTH-1:0] data_in;
    output logic [DATA_WIDTH-1:0] data_out;
);

    // sub_bytes
    // row shift
    // mix column
    // add key
    
endmodule